module IsNeg(input[15:0] in, output out);
  // your code here
 Or g1(in[15],1'b0,out);

endmodule
